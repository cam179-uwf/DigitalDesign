LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY bcd_10bit_decoder IS
	PORT (
		A,B,C,D				: IN STD_LOGIC;
		E,F,G,H,L,M,N,O,P,Q	: OUT STD_LOGIC;
		CLOCK: OUT STD_LOGIC
		);
END bcd_10bit_decoder;

ARCHITECTURE behaviour OF bcd_10bit_decoder IS
BEGIN
	Q <= NOT A AND NOT B AND NOT C AND NOT D;
	P <= NOT A AND NOT B AND NOT C AND D;
	O <= NOT A AND NOT B AND C AND NOT D;
	N <= NOT A AND NOT B AND C AND D;
	M <= NOT A AND B AND NOT C AND NOT D;
	L <= NOT A AND B AND NOT C AND D;
	H <= NOT A AND B AND C AND NOT D;
	G <= NOT A AND B AND C AND D;
	F <= A AND NOT B AND NOT C AND NOT D;
	E <= A AND NOT B AND NOT C AND D;
END behaviour;